library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pipeline is
 Port (
   clk : in std_logic;
   reset : in std_logic
   );
end pipeline;

architecture arch of pipeline is
begin

end arch;
